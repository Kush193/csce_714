//=====================================================================
// Project: 4 core MESI cache design
// File Name: read_miss_icache.sv
// Description: Test for back to back reads in same address in D-Cache
// Designers: Pranit, Aditya, Kushagra
//=====================================================================

class random_read_write_all_proc extends base_test;

    //component macro
    `uvm_component_utils(random_read_write_all_proc)

    //Constructor
    function new(string name, uvm_component parent);
        super.new(name, parent);
    endfunction : new

    //UVM build phase
    function void build_phase(uvm_phase phase);
        uvm_config_wrapper::set(this, "tb.vsequencer.run_phase", "default_sequence", random_read_write_all_proc_seq::type_id::get());
        super.build_phase(phase);
    endfunction : build_phase

    //UVM run phase()
    task run_phase(uvm_phase phase);
        `uvm_info(get_type_name(), "Executing random_read_write_all_proc test" , UVM_LOW)
    endtask: run_phase

endclass : random_read_write_all_proc


// Sequence for a read-miss on D-cache
class random_read_write_all_proc_seq extends base_vseq;
    //object macro
    `uvm_object_utils(random_read_write_all_proc_seq)
	bit [`ADDR_WID_LV1-1 : 0] addr;
    cpu_transaction_c trans;

    //constructor
    function new (string name="random_read_write_all_proc_seq");
        super.new(name);
    endfunction : new

    virtual task body();
        //trans.randomize();
        repeat(100) begin
        for(int i =0; i<4; i++)begin
            `uvm_do_on_with(trans, p_sequencer.cpu_seqr[i], {request_type == WRITE_REQ; access_cache_type == DCACHE_ACC;})
            addr = trans.address;
            `uvm_do_on_with(trans, p_sequencer.cpu_seqr[i], {request_type == READ_REQ; access_cache_type == DCACHE_ACC; address == addr;})

        end
        end
		
	endtask

endclass : random_read_write_all_proc_seq
